magic
tech gf180mcuD
magscale 1 5
timestamp 1700370116
<< obsm1 >>
rect 672 1538 279328 174078
<< metal2 >>
rect 139888 0 139944 400
<< obsm2 >>
rect 854 430 279258 174067
rect 854 400 139858 430
rect 139974 400 279258 430
<< metal3 >>
rect 279600 170240 280000 170296
rect 0 163184 400 163240
rect 279600 159264 280000 159320
rect 279600 148288 280000 148344
rect 0 138096 400 138152
rect 279600 137312 280000 137368
rect 279600 126336 280000 126392
rect 279600 115360 280000 115416
rect 0 113008 400 113064
rect 279600 104384 280000 104440
rect 279600 93408 280000 93464
rect 0 87920 400 87976
rect 279600 82432 280000 82488
rect 279600 71456 280000 71512
rect 0 62832 400 62888
rect 279600 60480 280000 60536
rect 279600 49504 280000 49560
rect 279600 38528 280000 38584
rect 0 37744 400 37800
rect 279600 27552 280000 27608
rect 279600 16576 280000 16632
rect 0 12656 400 12712
rect 279600 5600 280000 5656
<< obsm3 >>
rect 400 170326 279600 174062
rect 400 170210 279570 170326
rect 400 163270 279600 170210
rect 430 163154 279600 163270
rect 400 159350 279600 163154
rect 400 159234 279570 159350
rect 400 148374 279600 159234
rect 400 148258 279570 148374
rect 400 138182 279600 148258
rect 430 138066 279600 138182
rect 400 137398 279600 138066
rect 400 137282 279570 137398
rect 400 126422 279600 137282
rect 400 126306 279570 126422
rect 400 115446 279600 126306
rect 400 115330 279570 115446
rect 400 113094 279600 115330
rect 430 112978 279600 113094
rect 400 104470 279600 112978
rect 400 104354 279570 104470
rect 400 93494 279600 104354
rect 400 93378 279570 93494
rect 400 88006 279600 93378
rect 430 87890 279600 88006
rect 400 82518 279600 87890
rect 400 82402 279570 82518
rect 400 71542 279600 82402
rect 400 71426 279570 71542
rect 400 62918 279600 71426
rect 430 62802 279600 62918
rect 400 60566 279600 62802
rect 400 60450 279570 60566
rect 400 49590 279600 60450
rect 400 49474 279570 49590
rect 400 38614 279600 49474
rect 400 38498 279570 38614
rect 400 37830 279600 38498
rect 430 37714 279600 37830
rect 400 27638 279600 37714
rect 400 27522 279570 27638
rect 400 16662 279600 27522
rect 400 16546 279570 16662
rect 400 12742 279600 16546
rect 430 12626 279600 12742
rect 400 5686 279600 12626
rect 400 5570 279570 5686
rect 400 1554 279600 5570
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< obsm4 >>
rect 278614 77289 278674 104151
rect 278894 77289 279090 104151
<< labels >>
rlabel metal3 s 279600 5600 280000 5656 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 62832 400 62888 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 37744 400 37800 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 12656 400 12712 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 279600 27552 280000 27608 6 io_in[1]
port 5 nsew signal input
rlabel metal3 s 279600 49504 280000 49560 6 io_in[2]
port 6 nsew signal input
rlabel metal3 s 279600 71456 280000 71512 6 io_in[3]
port 7 nsew signal input
rlabel metal3 s 279600 93408 280000 93464 6 io_in[4]
port 8 nsew signal input
rlabel metal3 s 279600 115360 280000 115416 6 io_in[5]
port 9 nsew signal input
rlabel metal3 s 279600 137312 280000 137368 6 io_in[6]
port 10 nsew signal input
rlabel metal3 s 279600 159264 280000 159320 6 io_in[7]
port 11 nsew signal input
rlabel metal3 s 0 163184 400 163240 6 io_in[8]
port 12 nsew signal input
rlabel metal3 s 0 113008 400 113064 6 io_in[9]
port 13 nsew signal input
rlabel metal3 s 279600 16576 280000 16632 6 io_out[0]
port 14 nsew signal output
rlabel metal3 s 279600 38528 280000 38584 6 io_out[1]
port 15 nsew signal output
rlabel metal3 s 279600 60480 280000 60536 6 io_out[2]
port 16 nsew signal output
rlabel metal3 s 279600 82432 280000 82488 6 io_out[3]
port 17 nsew signal output
rlabel metal3 s 279600 104384 280000 104440 6 io_out[4]
port 18 nsew signal output
rlabel metal3 s 279600 126336 280000 126392 6 io_out[5]
port 19 nsew signal output
rlabel metal3 s 279600 148288 280000 148344 6 io_out[6]
port 20 nsew signal output
rlabel metal3 s 279600 170240 280000 170296 6 io_out[7]
port 21 nsew signal output
rlabel metal3 s 0 138096 400 138152 6 io_out[8]
port 22 nsew signal output
rlabel metal3 s 0 87920 400 87976 6 io_out[9]
port 23 nsew signal output
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 24 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 25 nsew ground bidirectional
rlabel metal2 s 139888 0 139944 400 6 wb_clk_i
port 26 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15279720
string GDS_FILE /root/work/caravel_user_project/openlane/ADC_LogiCompilation/runs/23_11_18_23_57/results/signoff/ADC_LogiCompilation.magic.gds
string GDS_START 230492
<< end >>

