magic
tech gf180mcuD
magscale 1 5
timestamp 1700369006
<< obsm1 >>
rect 672 1538 279328 174078
<< metal2 >>
rect 139888 0 139944 400
<< obsm2 >>
rect 854 430 279314 174067
rect 854 400 139858 430
rect 139974 400 279314 430
<< metal3 >>
rect 0 170912 400 170968
rect 279600 170240 280000 170296
rect 0 162176 400 162232
rect 279600 159264 280000 159320
rect 0 153440 400 153496
rect 279600 148288 280000 148344
rect 0 144704 400 144760
rect 279600 137312 280000 137368
rect 0 135968 400 136024
rect 0 127232 400 127288
rect 279600 126336 280000 126392
rect 0 118496 400 118552
rect 279600 115360 280000 115416
rect 0 109760 400 109816
rect 279600 104384 280000 104440
rect 0 101024 400 101080
rect 279600 93408 280000 93464
rect 0 92288 400 92344
rect 0 83552 400 83608
rect 279600 82432 280000 82488
rect 0 74816 400 74872
rect 279600 71456 280000 71512
rect 0 66080 400 66136
rect 279600 60480 280000 60536
rect 0 57344 400 57400
rect 279600 49504 280000 49560
rect 0 48608 400 48664
rect 0 39872 400 39928
rect 279600 38528 280000 38584
rect 0 31136 400 31192
rect 279600 27552 280000 27608
rect 0 22400 400 22456
rect 279600 16576 280000 16632
rect 0 13664 400 13720
rect 279600 5600 280000 5656
rect 0 4928 400 4984
<< obsm3 >>
rect 400 170998 279650 174062
rect 430 170882 279650 170998
rect 400 170326 279650 170882
rect 400 170210 279570 170326
rect 400 162262 279650 170210
rect 430 162146 279650 162262
rect 400 159350 279650 162146
rect 400 159234 279570 159350
rect 400 153526 279650 159234
rect 430 153410 279650 153526
rect 400 148374 279650 153410
rect 400 148258 279570 148374
rect 400 144790 279650 148258
rect 430 144674 279650 144790
rect 400 137398 279650 144674
rect 400 137282 279570 137398
rect 400 136054 279650 137282
rect 430 135938 279650 136054
rect 400 127318 279650 135938
rect 430 127202 279650 127318
rect 400 126422 279650 127202
rect 400 126306 279570 126422
rect 400 118582 279650 126306
rect 430 118466 279650 118582
rect 400 115446 279650 118466
rect 400 115330 279570 115446
rect 400 109846 279650 115330
rect 430 109730 279650 109846
rect 400 104470 279650 109730
rect 400 104354 279570 104470
rect 400 101110 279650 104354
rect 430 100994 279650 101110
rect 400 93494 279650 100994
rect 400 93378 279570 93494
rect 400 92374 279650 93378
rect 430 92258 279650 92374
rect 400 83638 279650 92258
rect 430 83522 279650 83638
rect 400 82518 279650 83522
rect 400 82402 279570 82518
rect 400 74902 279650 82402
rect 430 74786 279650 74902
rect 400 71542 279650 74786
rect 400 71426 279570 71542
rect 400 66166 279650 71426
rect 430 66050 279650 66166
rect 400 60566 279650 66050
rect 400 60450 279570 60566
rect 400 57430 279650 60450
rect 430 57314 279650 57430
rect 400 49590 279650 57314
rect 400 49474 279570 49590
rect 400 48694 279650 49474
rect 430 48578 279650 48694
rect 400 39958 279650 48578
rect 430 39842 279650 39958
rect 400 38614 279650 39842
rect 400 38498 279570 38614
rect 400 31222 279650 38498
rect 430 31106 279650 31222
rect 400 27638 279650 31106
rect 400 27522 279570 27638
rect 400 22486 279650 27522
rect 430 22370 279650 22486
rect 400 16662 279650 22370
rect 400 16546 279570 16662
rect 400 13750 279650 16546
rect 430 13634 279650 13750
rect 400 5686 279650 13634
rect 400 5570 279570 5686
rect 400 5014 279650 5570
rect 430 4898 279650 5014
rect 400 1554 279650 4898
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< obsm4 >>
rect 277998 39713 278474 125655
<< labels >>
rlabel metal3 s 0 162176 400 162232 6 BN[0]
port 1 nsew signal output
rlabel metal3 s 0 144704 400 144760 6 BN[1]
port 2 nsew signal output
rlabel metal3 s 0 127232 400 127288 6 BN[2]
port 3 nsew signal output
rlabel metal3 s 0 109760 400 109816 6 BN[3]
port 4 nsew signal output
rlabel metal3 s 0 92288 400 92344 6 BN[4]
port 5 nsew signal output
rlabel metal3 s 0 74816 400 74872 6 BN[5]
port 6 nsew signal output
rlabel metal3 s 0 57344 400 57400 6 BN[6]
port 7 nsew signal output
rlabel metal3 s 0 39872 400 39928 6 BN[7]
port 8 nsew signal output
rlabel metal3 s 0 22400 400 22456 6 BN[8]
port 9 nsew signal output
rlabel metal3 s 0 4928 400 4984 6 BN[9]
port 10 nsew signal output
rlabel metal3 s 0 170912 400 170968 6 B[0]
port 11 nsew signal output
rlabel metal3 s 0 153440 400 153496 6 B[1]
port 12 nsew signal output
rlabel metal3 s 0 135968 400 136024 6 B[2]
port 13 nsew signal output
rlabel metal3 s 0 118496 400 118552 6 B[3]
port 14 nsew signal output
rlabel metal3 s 0 101024 400 101080 6 B[4]
port 15 nsew signal output
rlabel metal3 s 0 83552 400 83608 6 B[5]
port 16 nsew signal output
rlabel metal3 s 0 66080 400 66136 6 B[6]
port 17 nsew signal output
rlabel metal3 s 0 48608 400 48664 6 B[7]
port 18 nsew signal output
rlabel metal3 s 0 31136 400 31192 6 B[8]
port 19 nsew signal output
rlabel metal3 s 0 13664 400 13720 6 B[9]
port 20 nsew signal output
rlabel metal3 s 279600 16576 280000 16632 6 CompN[0]
port 21 nsew signal input
rlabel metal3 s 279600 49504 280000 49560 6 CompN[1]
port 22 nsew signal input
rlabel metal3 s 279600 82432 280000 82488 6 CompN[2]
port 23 nsew signal input
rlabel metal3 s 279600 104384 280000 104440 6 CompN[3]
port 24 nsew signal input
rlabel metal3 s 279600 126336 280000 126392 6 CompN[4]
port 25 nsew signal input
rlabel metal3 s 279600 148288 280000 148344 6 CompN[5]
port 26 nsew signal input
rlabel metal3 s 279600 170240 280000 170296 6 CompN[6]
port 27 nsew signal input
rlabel metal3 s 279600 5600 280000 5656 6 Comp[0]
port 28 nsew signal input
rlabel metal3 s 279600 38528 280000 38584 6 Comp[1]
port 29 nsew signal input
rlabel metal3 s 279600 71456 280000 71512 6 Comp[2]
port 30 nsew signal input
rlabel metal3 s 279600 93408 280000 93464 6 Comp[3]
port 31 nsew signal input
rlabel metal3 s 279600 115360 280000 115416 6 Comp[4]
port 32 nsew signal input
rlabel metal3 s 279600 137312 280000 137368 6 Comp[5]
port 33 nsew signal input
rlabel metal3 s 279600 159264 280000 159320 6 Comp[6]
port 34 nsew signal input
rlabel metal3 s 279600 27552 280000 27608 6 Samp
port 35 nsew signal input
rlabel metal2 s 139888 0 139944 400 6 clk
port 36 nsew signal input
rlabel metal3 s 279600 60480 280000 60536 6 eoc
port 37 nsew signal output
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 38 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 39 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 39 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15123656
string GDS_FILE /root/work/caravel_user_project/openlane/ADC_Flash_Logic/runs/23_11_18_23_38/results/signoff/ADC_Flash_Logic.magic.gds
string GDS_START 170764
<< end >>

