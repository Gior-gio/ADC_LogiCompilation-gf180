VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ADC_LogiCompilation
  CLASS BLOCK ;
  FOREIGN ADC_LogiCompilation ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 56.000 2800.000 56.560 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.555000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 628.320 4.000 628.880 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.612000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 377.440 4.000 378.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.612000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.560 4.000 127.120 ;
    END
  END io_in[12]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 275.520 2800.000 276.080 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 495.040 2800.000 495.600 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 714.560 2800.000 715.120 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 934.080 2800.000 934.640 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1153.600 2800.000 1154.160 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1373.120 2800.000 1373.680 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1592.640 2800.000 1593.200 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1631.840 4.000 1632.400 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1130.080 4.000 1130.640 ;
    END
  END io_in[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 165.760 2800.000 166.320 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 385.280 2800.000 385.840 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 604.800 2800.000 605.360 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 824.320 2800.000 824.880 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1043.840 2800.000 1044.400 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1263.360 2800.000 1263.920 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1482.880 2800.000 1483.440 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1702.400 2800.000 1702.960 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1380.960 4.000 1381.520 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 879.200 4.000 879.760 ;
    END
  END io_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 1740.780 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 1740.780 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1398.880 0.000 1399.440 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 2793.280 1740.780 ;
      LAYER Metal2 ;
        RECT 8.540 4.300 2792.580 1740.670 ;
        RECT 8.540 4.000 1398.580 4.300 ;
        RECT 1399.740 4.000 2792.580 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1703.260 2796.000 1740.620 ;
        RECT 4.000 1702.100 2795.700 1703.260 ;
        RECT 4.000 1632.700 2796.000 1702.100 ;
        RECT 4.300 1631.540 2796.000 1632.700 ;
        RECT 4.000 1593.500 2796.000 1631.540 ;
        RECT 4.000 1592.340 2795.700 1593.500 ;
        RECT 4.000 1483.740 2796.000 1592.340 ;
        RECT 4.000 1482.580 2795.700 1483.740 ;
        RECT 4.000 1381.820 2796.000 1482.580 ;
        RECT 4.300 1380.660 2796.000 1381.820 ;
        RECT 4.000 1373.980 2796.000 1380.660 ;
        RECT 4.000 1372.820 2795.700 1373.980 ;
        RECT 4.000 1264.220 2796.000 1372.820 ;
        RECT 4.000 1263.060 2795.700 1264.220 ;
        RECT 4.000 1154.460 2796.000 1263.060 ;
        RECT 4.000 1153.300 2795.700 1154.460 ;
        RECT 4.000 1130.940 2796.000 1153.300 ;
        RECT 4.300 1129.780 2796.000 1130.940 ;
        RECT 4.000 1044.700 2796.000 1129.780 ;
        RECT 4.000 1043.540 2795.700 1044.700 ;
        RECT 4.000 934.940 2796.000 1043.540 ;
        RECT 4.000 933.780 2795.700 934.940 ;
        RECT 4.000 880.060 2796.000 933.780 ;
        RECT 4.300 878.900 2796.000 880.060 ;
        RECT 4.000 825.180 2796.000 878.900 ;
        RECT 4.000 824.020 2795.700 825.180 ;
        RECT 4.000 715.420 2796.000 824.020 ;
        RECT 4.000 714.260 2795.700 715.420 ;
        RECT 4.000 629.180 2796.000 714.260 ;
        RECT 4.300 628.020 2796.000 629.180 ;
        RECT 4.000 605.660 2796.000 628.020 ;
        RECT 4.000 604.500 2795.700 605.660 ;
        RECT 4.000 495.900 2796.000 604.500 ;
        RECT 4.000 494.740 2795.700 495.900 ;
        RECT 4.000 386.140 2796.000 494.740 ;
        RECT 4.000 384.980 2795.700 386.140 ;
        RECT 4.000 378.300 2796.000 384.980 ;
        RECT 4.300 377.140 2796.000 378.300 ;
        RECT 4.000 276.380 2796.000 377.140 ;
        RECT 4.000 275.220 2795.700 276.380 ;
        RECT 4.000 166.620 2796.000 275.220 ;
        RECT 4.000 165.460 2795.700 166.620 ;
        RECT 4.000 127.420 2796.000 165.460 ;
        RECT 4.300 126.260 2796.000 127.420 ;
        RECT 4.000 56.860 2796.000 126.260 ;
        RECT 4.000 55.700 2795.700 56.860 ;
        RECT 4.000 15.540 2796.000 55.700 ;
      LAYER Metal4 ;
        RECT 2786.140 772.890 2786.740 1041.510 ;
        RECT 2788.940 772.890 2790.900 1041.510 ;
  END
END ADC_LogiCompilation
END LIBRARY

