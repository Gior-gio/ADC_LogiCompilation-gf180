VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ADC_Flash_Logic
  CLASS BLOCK ;
  FOREIGN ADC_Flash_Logic ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN BN[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1621.760 4.000 1622.320 ;
    END
  END BN[0]
  PIN BN[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1447.040 4.000 1447.600 ;
    END
  END BN[1]
  PIN BN[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1272.320 4.000 1272.880 ;
    END
  END BN[2]
  PIN BN[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1097.600 4.000 1098.160 ;
    END
  END BN[3]
  PIN BN[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 922.880 4.000 923.440 ;
    END
  END BN[4]
  PIN BN[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 748.160 4.000 748.720 ;
    END
  END BN[5]
  PIN BN[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 573.440 4.000 574.000 ;
    END
  END BN[6]
  PIN BN[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 398.720 4.000 399.280 ;
    END
  END BN[7]
  PIN BN[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.000 4.000 224.560 ;
    END
  END BN[8]
  PIN BN[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.280 4.000 49.840 ;
    END
  END BN[9]
  PIN B[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1709.120 4.000 1709.680 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1534.400 4.000 1534.960 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1359.680 4.000 1360.240 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1184.960 4.000 1185.520 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1010.240 4.000 1010.800 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 835.520 4.000 836.080 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 660.800 4.000 661.360 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 486.080 4.000 486.640 ;
    END
  END B[7]
  PIN B[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 311.360 4.000 311.920 ;
    END
  END B[8]
  PIN B[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 136.640 4.000 137.200 ;
    END
  END B[9]
  PIN CompN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 165.760 2800.000 166.320 ;
    END
  END CompN[0]
  PIN CompN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 495.040 2800.000 495.600 ;
    END
  END CompN[1]
  PIN CompN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 824.320 2800.000 824.880 ;
    END
  END CompN[2]
  PIN CompN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1043.840 2800.000 1044.400 ;
    END
  END CompN[3]
  PIN CompN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1263.360 2800.000 1263.920 ;
    END
  END CompN[4]
  PIN CompN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1482.880 2800.000 1483.440 ;
    END
  END CompN[5]
  PIN CompN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1702.400 2800.000 1702.960 ;
    END
  END CompN[6]
  PIN Comp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 56.000 2800.000 56.560 ;
    END
  END Comp[0]
  PIN Comp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 385.280 2800.000 385.840 ;
    END
  END Comp[1]
  PIN Comp[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 714.560 2800.000 715.120 ;
    END
  END Comp[2]
  PIN Comp[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 934.080 2800.000 934.640 ;
    END
  END Comp[3]
  PIN Comp[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1153.600 2800.000 1154.160 ;
    END
  END Comp[4]
  PIN Comp[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1373.120 2800.000 1373.680 ;
    END
  END Comp[5]
  PIN Comp[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1592.640 2800.000 1593.200 ;
    END
  END Comp[6]
  PIN Samp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 275.520 2800.000 276.080 ;
    END
  END Samp
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.555000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1398.880 0.000 1399.440 4.000 ;
    END
  END clk
  PIN eoc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 604.800 2800.000 605.360 ;
    END
  END eoc
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 1740.780 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 1740.780 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 2793.280 1740.780 ;
      LAYER Metal2 ;
        RECT 8.540 4.300 2793.140 1740.670 ;
        RECT 8.540 4.000 1398.580 4.300 ;
        RECT 1399.740 4.000 2793.140 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1709.980 2796.500 1740.620 ;
        RECT 4.300 1708.820 2796.500 1709.980 ;
        RECT 4.000 1703.260 2796.500 1708.820 ;
        RECT 4.000 1702.100 2795.700 1703.260 ;
        RECT 4.000 1622.620 2796.500 1702.100 ;
        RECT 4.300 1621.460 2796.500 1622.620 ;
        RECT 4.000 1593.500 2796.500 1621.460 ;
        RECT 4.000 1592.340 2795.700 1593.500 ;
        RECT 4.000 1535.260 2796.500 1592.340 ;
        RECT 4.300 1534.100 2796.500 1535.260 ;
        RECT 4.000 1483.740 2796.500 1534.100 ;
        RECT 4.000 1482.580 2795.700 1483.740 ;
        RECT 4.000 1447.900 2796.500 1482.580 ;
        RECT 4.300 1446.740 2796.500 1447.900 ;
        RECT 4.000 1373.980 2796.500 1446.740 ;
        RECT 4.000 1372.820 2795.700 1373.980 ;
        RECT 4.000 1360.540 2796.500 1372.820 ;
        RECT 4.300 1359.380 2796.500 1360.540 ;
        RECT 4.000 1273.180 2796.500 1359.380 ;
        RECT 4.300 1272.020 2796.500 1273.180 ;
        RECT 4.000 1264.220 2796.500 1272.020 ;
        RECT 4.000 1263.060 2795.700 1264.220 ;
        RECT 4.000 1185.820 2796.500 1263.060 ;
        RECT 4.300 1184.660 2796.500 1185.820 ;
        RECT 4.000 1154.460 2796.500 1184.660 ;
        RECT 4.000 1153.300 2795.700 1154.460 ;
        RECT 4.000 1098.460 2796.500 1153.300 ;
        RECT 4.300 1097.300 2796.500 1098.460 ;
        RECT 4.000 1044.700 2796.500 1097.300 ;
        RECT 4.000 1043.540 2795.700 1044.700 ;
        RECT 4.000 1011.100 2796.500 1043.540 ;
        RECT 4.300 1009.940 2796.500 1011.100 ;
        RECT 4.000 934.940 2796.500 1009.940 ;
        RECT 4.000 933.780 2795.700 934.940 ;
        RECT 4.000 923.740 2796.500 933.780 ;
        RECT 4.300 922.580 2796.500 923.740 ;
        RECT 4.000 836.380 2796.500 922.580 ;
        RECT 4.300 835.220 2796.500 836.380 ;
        RECT 4.000 825.180 2796.500 835.220 ;
        RECT 4.000 824.020 2795.700 825.180 ;
        RECT 4.000 749.020 2796.500 824.020 ;
        RECT 4.300 747.860 2796.500 749.020 ;
        RECT 4.000 715.420 2796.500 747.860 ;
        RECT 4.000 714.260 2795.700 715.420 ;
        RECT 4.000 661.660 2796.500 714.260 ;
        RECT 4.300 660.500 2796.500 661.660 ;
        RECT 4.000 605.660 2796.500 660.500 ;
        RECT 4.000 604.500 2795.700 605.660 ;
        RECT 4.000 574.300 2796.500 604.500 ;
        RECT 4.300 573.140 2796.500 574.300 ;
        RECT 4.000 495.900 2796.500 573.140 ;
        RECT 4.000 494.740 2795.700 495.900 ;
        RECT 4.000 486.940 2796.500 494.740 ;
        RECT 4.300 485.780 2796.500 486.940 ;
        RECT 4.000 399.580 2796.500 485.780 ;
        RECT 4.300 398.420 2796.500 399.580 ;
        RECT 4.000 386.140 2796.500 398.420 ;
        RECT 4.000 384.980 2795.700 386.140 ;
        RECT 4.000 312.220 2796.500 384.980 ;
        RECT 4.300 311.060 2796.500 312.220 ;
        RECT 4.000 276.380 2796.500 311.060 ;
        RECT 4.000 275.220 2795.700 276.380 ;
        RECT 4.000 224.860 2796.500 275.220 ;
        RECT 4.300 223.700 2796.500 224.860 ;
        RECT 4.000 166.620 2796.500 223.700 ;
        RECT 4.000 165.460 2795.700 166.620 ;
        RECT 4.000 137.500 2796.500 165.460 ;
        RECT 4.300 136.340 2796.500 137.500 ;
        RECT 4.000 56.860 2796.500 136.340 ;
        RECT 4.000 55.700 2795.700 56.860 ;
        RECT 4.000 50.140 2796.500 55.700 ;
        RECT 4.300 48.980 2796.500 50.140 ;
        RECT 4.000 15.540 2796.500 48.980 ;
      LAYER Metal4 ;
        RECT 2779.980 397.130 2784.740 1256.550 ;
  END
END ADC_Flash_Logic
END LIBRARY

